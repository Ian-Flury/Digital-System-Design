library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.all;


entity lcd_ctrl_top is
    port(
        clock_50M   : in std_logic;
        KEY3        : in std_logic
    );
end lcd_ctrl_top;

architecture structural of lcd_ctrl_top is

begin

end structural;
