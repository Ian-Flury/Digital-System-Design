library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.all;

entity lcd_ctrl is

end lcd_ctrl;


architecture rtl of lcd_ctrl is 

begin

end rtl;